module csa(
    input [7:0]input_1,
    input [7:0]input_2,
    output [7:0]add_out,
    output [7:0]add_overflow
    );
endmodule